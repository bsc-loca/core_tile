
module sim_top;
    import sargantana_hpdc_pkg::*, drac_pkg::*;

    logic tb_clk, tb_rstn;

    // *** Clock & Reset drivers ***

    initial begin
        tb_clk = 1'b0;
        tb_rstn = 1'b0;
        #5 tb_rstn = 1'b1;
    end

    always #1 tb_clk = ~tb_clk;

    // *** DUT ***


    // Bootrom wires
    logic [23:0] brom_req_address;
    logic brom_req_valid;
    logic brom_ready;
    logic [127:0] brom_resp_data;
    logic brom_resp_valid;

    // icache wires
    logic icache_l1_request_valid;
    logic icache_l2_response_valid;
    logic [drac_pkg::PHY_ADDR_SIZE-1:0] icache_l1_request_paddr;
    logic [sargantana_icache_pkg::FETCH_WIDHT-1:0] icache_l2_response_data;

    logic dut_icache_req_valid;
    logic dut_icache_resp_valid;
    logic [drac_pkg::PHY_ADDR_SIZE-1:0] dut_icache_request_paddr;
    logic [sargantana_icache_pkg::FETCH_WIDHT-1:0] dut_icache_response_data;

    assign dut_icache_response_data = brom_resp_valid ? brom_resp_data : icache_l2_response_data;
    assign dut_icache_response_valid = brom_resp_valid | icache_l2_response_valid;
    assign icache_l1_request_paddr = dut_icache_request_paddr;
    assign icache_l1_request_valid = dut_icache_req_valid;

    //      Miss read interface
    logic                          mem_req_miss_read_ready;
    logic                          mem_req_miss_read_valid;
    hpdcache_mem_req_t             mem_req_miss_read;

    logic                          mem_resp_miss_read_ready;
    logic                          mem_resp_miss_read_valid;
    hpdcache_mem_resp_r_t          mem_resp_miss_read;

    //      Write-buffer write interface
    logic                          mem_req_wbuf_write_ready;
    logic                          mem_req_wbuf_write_valid;
    hpdcache_mem_req_t             mem_req_wbuf_write;

    logic                          mem_req_wbuf_write_data_ready;
    logic                          mem_req_wbuf_write_data_valid;
    hpdcache_mem_req_w_t           mem_req_wbuf_write_data;

    logic                          mem_resp_wbuf_write_ready;
    logic                          mem_resp_wbuf_write_valid;
    hpdcache_mem_resp_w_t          mem_resp_wbuf_write;

    //      Uncached read interface
    logic                          mem_req_uc_read_ready;
    logic                          mem_req_uc_read_valid;
    hpdcache_mem_req_t             mem_req_uc_read;

    logic                          mem_resp_uc_read_ready;
    logic                          mem_resp_uc_read_valid;
    hpdcache_mem_resp_r_t          mem_resp_uc_read;

    //      Uncached write interface
    logic                          mem_req_uc_write_ready;
    logic                          mem_req_uc_write_valid;
    hpdcache_mem_req_t             mem_req_uc_write;

    logic                          mem_req_uc_write_data_ready;
    logic                          mem_req_uc_write_data_valid;
    hpdcache_mem_req_w_t           mem_req_uc_write_data;

    logic                          mem_resp_uc_write_ready;
    logic                          mem_resp_uc_write_valid;
    hpdcache_mem_resp_w_t          mem_resp_uc_write;

    // Debug Module Interface

    // DM -> Core
    debug_contr_in_t debug_contr_dm_to_core;
    debug_reg_in_t   debug_reg_dm_to_core;

    // Core -> DM
    debug_contr_out_t debug_contr_core_to_dm;
    debug_reg_out_t   debug_reg_core_to_dm;

    logic dut_rstn, debug_reset;

    assign dut_rstn = ~(~tb_rstn | debug_reset);

    top_tile DUT(
        .clk_i(tb_clk),
        .rstn_i(dut_rstn),
        .soft_rstn_i(dut_rstn),
        .reset_addr_i({{{PHY_VIRT_MAX_ADDR_SIZE-16}{1'b0}}, 16'h0100}),
        .core_id_i(64'b0),

        // Bootrom ports
        .brom_req_address_o(brom_req_address),
        .brom_req_valid_o(brom_req_valid),

        // icache ports
        .io_mem_acquire_valid(dut_icache_req_valid),               
        .io_mem_acquire_bits_addr_block(dut_icache_request_paddr),   
        .io_mem_grant_valid(dut_icache_response_valid),         
        .io_mem_grant_bits_data(dut_icache_response_data),
        .io_mem_grant_inval(0),
        .io_mem_grant_inval_addr(0),

        // dmem ports

        // dMem miss-read interface
        .mem_req_miss_read_ready_i(mem_req_miss_read_ready),
        .mem_req_miss_read_valid_o(mem_req_miss_read_valid),
        .mem_req_miss_read_o(mem_req_miss_read),

        .mem_resp_miss_read_ready_o(mem_resp_miss_read_ready),
        .mem_resp_miss_read_valid_i(mem_resp_miss_read_valid),
        .mem_resp_miss_read_i(mem_resp_miss_read),

        // dMem writeback interface
        .mem_req_wbuf_write_ready_i(mem_req_wbuf_write_ready),
        .mem_req_wbuf_write_valid_o(mem_req_wbuf_write_valid),
        .mem_req_wbuf_write_o(mem_req_wbuf_write),

        .mem_req_wbuf_write_data_ready_i(mem_req_wbuf_write_data_ready),
        .mem_req_wbuf_write_data_valid_o(mem_req_wbuf_write_data_valid),
        .mem_req_wbuf_write_data_o(mem_req_wbuf_write_data),

        .mem_resp_wbuf_write_ready_o(mem_resp_wbuf_write_ready),
        .mem_resp_wbuf_write_valid_i(mem_resp_wbuf_write_valid),
        .mem_resp_wbuf_write_i(mem_resp_wbuf_write),

        // dMem uncacheable write interface
        .mem_req_uc_write_ready_i(mem_req_uc_write_ready),
        .mem_req_uc_write_valid_o(mem_req_uc_write_valid),
        .mem_req_uc_write_o(mem_req_uc_write),

        .mem_req_uc_write_data_ready_i(mem_req_uc_write_data_ready),
        .mem_req_uc_write_data_valid_o(mem_req_uc_write_data_valid),
        .mem_req_uc_write_data_o(mem_req_uc_write_data),

        .mem_resp_uc_write_ready_o(mem_resp_uc_write_ready),
        .mem_resp_uc_write_valid_i(mem_resp_uc_write_valid),
        .mem_resp_uc_write_i(mem_resp_uc_write),

        // dMem uncacheable read interface
        .mem_req_uc_read_ready_i(mem_req_uc_read_ready),
        .mem_req_uc_read_valid_o(mem_req_uc_read_valid),
        .mem_req_uc_read_o(mem_req_uc_read),

        .mem_resp_uc_read_ready_o(mem_resp_uc_read_ready),
        .mem_resp_uc_read_valid_i(mem_resp_uc_read_valid),
        .mem_resp_uc_read_i(mem_resp_uc_read),

        // Unused ports
        
        .debug_contr_i(debug_contr_dm_to_core),
        .debug_reg_i(debug_reg_dm_to_core),
        .debug_contr_o(debug_contr_core_to_dm),
        .debug_reg_o(debug_reg_core_to_dm),

        .time_i(64'd0),
        .irq_i(1'b0),
        .soft_irq_i(1'b0),
        .time_irq_i(1'b0),
        .io_core_pmu_l2_hit_i()
    );

    // *** Bootrom ***

    bootrom_behav brom(
        .clk(tb_clk),
        .rstn(tb_rstn),
        .brom_req_address_i(brom_req_address),
        .brom_req_valid_i(brom_req_valid),
        .brom_ready_o(brom_ready),
        .brom_resp_data_o(brom_resp_data),
        .brom_resp_valid_o(brom_resp_valid)
    );

    // *** L2 / Main Memory ***

    l2_behav #(
        .DATA_CACHE_LINE_SIZE(drac_pkg::DCACHE_BUS_WIDTH),
        .INST_CACHE_LINE_SIZE(sargantana_icache_pkg::SET_WIDHT)
    ) l2_inst (
        .clk_i(tb_clk),
        .rstn_i(tb_rstn),

        // *** Instruction Cache Interface ***

        .ic_addr_i(icache_l1_request_paddr),
        .ic_valid_i(icache_l1_request_valid),
        .ic_valid_o(icache_l2_response_valid),
        .ic_line_o(icache_l2_response_data),
	    .ic_seq_num_o(),

        // *** dCache Miss Read Interface ***

        .dc_mr_addr_i(mem_req_miss_read.mem_req_addr),
        .dc_mr_valid_i(mem_req_miss_read_valid),
        .dc_mr_ready_i(mem_resp_miss_read_ready),
        .dc_mr_tag_i(mem_req_miss_read.mem_req_id),
        .dc_mr_word_size_i(mem_req_miss_read.mem_req_size),
        .dc_mr_data_o(mem_resp_miss_read.mem_resp_r_data),
        .dc_mr_ready_o(mem_req_miss_read_ready),
        .dc_mr_valid_o(mem_resp_miss_read_valid),
        .dc_mr_tag_o(mem_resp_miss_read.mem_resp_r_id),
        .dc_mr_last_o(mem_resp_miss_read.mem_resp_r_last),

        // *** dCache Writeback Interface ***
        .dc_wb_req_ready_o(mem_req_wbuf_write_ready),
        .dc_wb_req_valid_i(mem_req_wbuf_write_valid),
        .dc_wb_req_addr_i(mem_req_wbuf_write.mem_req_addr),
        .dc_wb_req_len_i(mem_req_wbuf_write.mem_req_len),
        .dc_wb_req_size_i(mem_req_wbuf_write.mem_req_size),
        .dc_wb_req_id_i(mem_req_wbuf_write.mem_req_id),

        .dc_wb_req_data_ready_o(mem_req_wbuf_write_data_ready),
        .dc_wb_req_data_valid_i(mem_req_wbuf_write_data_valid),
        .dc_wb_req_data_i(mem_req_wbuf_write_data.mem_req_w_data),
        .dc_wb_req_be_i(mem_req_wbuf_write_data.mem_req_w_be),
        .dc_wb_req_last_i(mem_req_wbuf_write_data.mem_req_w_last),

        .dc_wb_resp_ready_i(mem_resp_wbuf_write_ready),
        .dc_wb_resp_valid_o(mem_resp_wbuf_write_valid),
        .dc_wb_resp_error_o(mem_resp_wbuf_write.mem_resp_w_error),
        .dc_wb_resp_id_o(mem_resp_wbuf_write.mem_resp_w_id),

        // *** dCache Uncacheable Writes Interface ***
        .dc_uc_wr_req_ready_o(mem_req_uc_write_ready),
        .dc_uc_wr_req_valid_i(mem_req_uc_write_valid),
        .dc_uc_wr_req_addr_i(mem_req_uc_write.mem_req_addr),
        .dc_uc_wr_req_len_i(mem_req_uc_write.mem_req_len),
        .dc_uc_wr_req_size_i(mem_req_uc_write.mem_req_size),
        .dc_uc_wr_req_id_i(mem_req_uc_write.mem_req_id),
        .dc_uc_wr_req_command_i(mem_req_uc_write.mem_req_command),
        .dc_uc_wr_req_atomic_i(mem_req_uc_write.mem_req_atomic),

        .dc_uc_wr_req_data_ready_o(mem_req_uc_write_data_ready),
        .dc_uc_wr_req_data_valid_i(mem_req_uc_write_data_valid),
        .dc_uc_wr_req_data_i(mem_req_uc_write_data.mem_req_w_data),
        .dc_uc_wr_req_be_i(mem_req_uc_write_data.mem_req_w_be),
        .dc_uc_wr_req_last_i(mem_req_uc_write_data.mem_req_w_last),

        .dc_uc_wr_resp_ready_i(mem_resp_uc_write_ready),
        .dc_uc_wr_resp_valid_o(mem_resp_uc_write_valid),
        .dc_uc_wr_resp_is_atomic_o(mem_resp_uc_write.mem_resp_w_is_atomic),
        .dc_uc_wr_resp_error_o(mem_resp_uc_write.mem_resp_w_error),
        .dc_uc_wr_resp_id_o(mem_resp_uc_write.mem_resp_w_id),

        // *** dCache Uncacheable Reads Interface ***
        .dc_uc_rd_req_ready_o(mem_req_uc_read_ready),
        .dc_uc_rd_req_valid_i(mem_req_uc_read_valid),
        .dc_uc_rd_req_addr_i(mem_req_uc_read.mem_req_addr),
        .dc_uc_rd_req_len_i(mem_req_uc_read.mem_req_len),
        .dc_uc_rd_req_size_i(mem_req_uc_read.mem_req_size),
        .dc_uc_rd_req_id_i(mem_req_uc_read.mem_req_id),
        .dc_uc_rd_req_command_i(mem_req_uc_read.mem_req_command),
        .dc_uc_rd_req_atomic_i(mem_req_uc_read.mem_req_atomic),

        .dc_uc_rd_valid_o(mem_resp_uc_read_valid),
        .dc_uc_rd_error_o(mem_resp_uc_read_error),
        .dc_uc_rd_id_o(mem_resp_uc_read.mem_resp_r_id),
        .dc_uc_rd_data_o(mem_resp_uc_read.mem_resp_r_data),
        .dc_uc_rd_last_o(mem_resp_uc_read.mem_resp_r_last),
        .dc_uc_rd_ready_i(mem_resp_uc_read_ready)
    );

    // Debug Module / JTAG

    logic tck, tms, tdi, tdo, trstn, tdo_driven, jtag_enable;

    SimJTAG #(
        .TICK_DELAY(0)
    ) JTAG_DPI (
        .clock(tb_clk),
        .reset(~tb_rstn),

        .enable(jtag_enable),
        .init_done(1),

        .jtag_TCK(tck),
        .jtag_TMS(tms),
        .jtag_TDI(tdi),
        .jtag_TRSTn(trstn),

        .jtag_TDO_data(tdo),
        .jtag_TDO_driven(tdo_driven),

        .exit()
    );

    logic                                       req_valid;
    logic                                       req_ready;
    logic [riscv_dm_pkg::DMI_ADDR_WIDTH-1:0]    req_addr;
    logic [riscv_dm_pkg::DMI_DATA_WIDTH-1:0]    req_data;
    logic [riscv_dm_pkg::DMI_OP_WIDTH-1:0]      req_op;
    logic                                       req_valid_cdc;
    logic                                       req_ready_cdc;
    logic [riscv_dm_pkg::DMI_ADDR_WIDTH-1:0]    req_addr_cdc;
    logic [riscv_dm_pkg::DMI_DATA_WIDTH-1:0]    req_data_cdc;
    logic [riscv_dm_pkg::DMI_OP_WIDTH-1:0]      req_op_cdc;

    logic                                       resp_valid;
    logic                                       resp_ready;
    logic [riscv_dm_pkg::DMI_DATA_WIDTH-1:0]    resp_data;
    logic [riscv_dm_pkg::DMI_OP_WIDTH-1:0]      resp_op;
    logic                                       resp_valid_cdc;
    logic                                       resp_ready_cdc;
    logic [riscv_dm_pkg::DMI_DATA_WIDTH-1:0]    resp_data_cdc;
    logic [riscv_dm_pkg::DMI_OP_WIDTH-1:0]      resp_op_cdc;

    riscv_dtm dtm(
        .tms_i(tms),
        .tck_i(tck),
        .trst_i(~trstn),
        .tdi_i(tdi),
        .tdo_o(tdo),
        .tdo_driven_o(tdo_driven),

        .req_valid_o(req_valid),
        .req_ready_i(req_ready),
        .req_addr_o(req_addr),
        .req_data_o(req_data),
        .req_op_o(req_op),

        .resp_valid_i(resp_valid_cdc),
        .resp_ready_o(resp_ready_cdc),
        .resp_data_i(resp_data_cdc),
        .resp_op_i(resp_op_cdc)
    );

    cdc_fifo_gray_clearable #(
        .WIDTH(riscv_dm_pkg::DMI_ADDR_WIDTH+riscv_dm_pkg::DMI_DATA_WIDTH+riscv_dm_pkg::DMI_OP_WIDTH)
    ) req_cdc_fifo (
        .src_rst_ni(trstn),
        .src_clk_i(tck),
        .src_clear_i(0),
        .src_clear_pending_o(),
        .src_data_i({req_addr, req_data, req_op}),
        .src_valid_i(req_valid),
        .src_ready_o(req_ready),

        .dst_rst_ni(tb_rstn),
        .dst_clk_i(tb_clk),
        .dst_clear_i(0),
        .dst_clear_pending_o(),
        .dst_data_o({req_addr_cdc, req_data_cdc, req_op_cdc}),
        .dst_valid_o(req_valid_cdc),
        .dst_ready_i(req_ready_cdc)
    );

    cdc_fifo_gray_clearable #(
        .WIDTH(riscv_dm_pkg::DMI_DATA_WIDTH+riscv_dm_pkg::DMI_OP_WIDTH)
    ) resp_cdc_fifo (
        .src_rst_ni(tb_rstn),
        .src_clk_i(tb_clk),
        .src_clear_i(0),
        .src_clear_pending_o(),
        .src_data_i({resp_data, resp_op}),
        .src_valid_i(resp_valid),
        .src_ready_o(resp_ready),

        .dst_rst_ni(trstn),
        .dst_clk_i(tck),
        .dst_clear_i(0),
        .dst_clear_pending_o(),
        .dst_data_o({resp_data_cdc, resp_op_cdc}),
        .dst_valid_o(resp_valid_cdc),
        .dst_ready_i(resp_ready_cdc)
    );

    logic halt_request, resume_request, halted, resumeack;

    riscv_dm dm(
        .clk_i(tb_clk),
        .rstn_i(tb_rstn),

        .req_valid_i(req_valid_cdc),
        .req_ready_o(req_ready_cdc),
        .req_addr_i(req_addr_cdc),
        .req_data_i(req_data_cdc),
        .req_op_i(req_op_cdc),

        .resp_valid_o(resp_valid),
        .resp_ready_i(resp_ready),
        .resp_data_o(resp_data),
        .resp_op_o(resp_op),

        .resume_request_o(debug_contr_dm_to_core.resume_req),
        .halt_request_o(debug_contr_dm_to_core.halt_req),
        .halt_on_reset_o(debug_contr_dm_to_core.halt_on_reset),
        .progbuf_run_req_o(debug_contr_dm_to_core.progbuf_req),
        .hart_reset_o(debug_reset),

        .resume_ack_i(debug_contr_core_to_dm.resume_ack),
        .halted_i(debug_contr_core_to_dm.halted),
        .running_i(debug_contr_core_to_dm.running),
        .havereset_i(0),
        .unavail_i(debug_contr_core_to_dm.unavail),
        .progbuf_run_ack_i(debug_contr_core_to_dm.progbuf_ack),
        .parked_i(debug_contr_core_to_dm.parked),

        .rnm_read_en_o(debug_reg_dm_to_core.rnm_read_en),       // Request reading the rename table
        .rnm_read_reg_o(debug_reg_dm_to_core.rnm_read_reg),     // Logical register for which the mapping is read
        .rnm_read_resp_i(debug_reg_core_to_dm.rnm_read_resp),   // Physical register mapped to the requested logical register

        .rf_en_o(debug_reg_dm_to_core.rf_en),                   // Read enable for the register file
        .rf_preg_o(debug_reg_dm_to_core.rf_preg),               // Target physical register in the register file
        .rf_rdata_i(debug_reg_core_to_dm.rf_rdata),             // Data read from the register file

        .rf_we_o(debug_reg_dm_to_core.rf_we),                   // Write enable for the register file
        .rf_wdata_o(debug_reg_dm_to_core.rf_wdata),             // Data to write to the register file
        //! @end


        // SRI interface for program buffer
        //! @virtualbus sri @dir in
        .sri_addr_i('0),     //! register interface address
        .sri_en_i('0),       //! register interface enable
        .sri_wdata_i('0),    //! register interface data to write
        .sri_we_i('0),       //! register interface write enable
        .sri_be_i('0),       //! register interface byte enable
        .sri_rdata_o(),    //! register interface read data
        .sri_error_o()     //! register interface error
    );

    // *** Testbench monitors ***

    logic [63:0] cycles, max_cycles, start_cycles;

    always @(posedge tb_clk, negedge tb_rstn) begin
        if (~tb_rstn) cycles <= 0;
        else cycles <= cycles + 1;
    end

    initial begin
        string dumpfile;
        start_cycles = 0;
        if ($test$plusargs("vcd")) begin
            $dumpfile("dump_file.vcd");
            if (!$value$plusargs("start-vcd-cycles=%d", start_cycles)) begin
                $dumpvars();
            end
        end
        if (!$value$plusargs("max-cycles=%d", max_cycles)) max_cycles = 0;
    end

    always @(posedge tb_clk) begin
        if (start_cycles > 0 && cycles == start_cycles) begin
            $dumpvars();
        end
    end

    always @(posedge tb_clk) begin
        if (max_cycles > 0 && cycles == max_cycles) begin
            $error("Test timeout");
            $finish;
        end
    end

    initial begin
        if ($test$plusargs("jtag")) begin
            jtag_enable = 1'b1;
        end else begin
            jtag_enable = 1'b0;
        end
    end

endmodule // veri_top
