//`default_nettype none
//`include "drac_pkg.sv"

/* -----------------------------------------------
 * Project Name   : DRAC
 * File           : mem_unit.v
 * Organization   : Barcelona Supercomputing Center
 * Author(s)      : Rubén Langarita
 * Email(s)       : ruben.langarita@bsc.es
 * -----------------------------------------------
 * Revision History
 *  Revision   | Author     | Description
 *  0.1        | Ruben. L   |
 *  0.2        | Victor. SP | Improve Doc. and pass tb
 *  0.3        | Arnau B.   | Modify to work with HPDC
 * -----------------------------------------------
 */
 
// Interface with Data Cache. Stores a Memory request until it finishes

module dcache_interface 
    import drac_pkg::*, hpdcache_pkg::*;
#(
    parameter drac_pkg::drac_cfg_t DracCfg     = drac_pkg::DracDefaultConfig
)(
    input  logic                clk_i,             // Clock
    input  logic                rstn_i,            // Negative Reset Signal

    // CPU Interface
    input  req_cpu_dcache_t     req_cpu_dcache_i,
    output resp_dcache_cpu_t    resp_dcache_cpu_o, // Dcache to CPU

    // dCache Interface
    input  logic dcache_ready_i,
    input  logic dcache_valid_i,
    output logic core_req_valid_o,
    output hpdcache_req_t req_dcache_o,
    output logic req_dcache_abort_o,
    output hpdcache_tag_t req_dcache_tag_o,
    output hpdcache_pma_t req_dcache_pma_o,
    input  hpdcache_rsp_t rsp_dcache_i,
    input logic wbuf_empty_i,

    // PMU
    output logic                dmem_is_store_o,
    output logic                dmem_is_load_o
);

logic io_address_space;

// The address is in the INPUT/OUTPUT space
assign io_address_space = (is_inside_IO_sections(DracCfg, req_cpu_dcache_i.data_rs1));

//-------------------------------------------------------------
// dCache Interface
//-------------------------------------------------------------

logic wait_resp_same_tag; // This signal identifies when the core must wait for
                          // the cache to process an old request with the same
                          // tag that's about to be used for the next request.

assign core_req_valid_o = req_cpu_dcache_i.valid & ~wait_resp_same_tag; 

// Memory Operation
always_comb begin
    case(req_cpu_dcache_i.instr_type)
        AMO_LRW,AMO_LRD:     req_dcache_o.op = HPDCACHE_REQ_AMO_LR;
        AMO_SCW,AMO_SCD:     req_dcache_o.op = HPDCACHE_REQ_AMO_SC;
        AMO_SWAPW,AMO_SWAPD: req_dcache_o.op = HPDCACHE_REQ_AMO_SWAP;
        AMO_ADDW,AMO_ADDD:   req_dcache_o.op = HPDCACHE_REQ_AMO_ADD;
        AMO_XORW,AMO_XORD:   req_dcache_o.op = HPDCACHE_REQ_AMO_XOR;
        AMO_ANDW,AMO_ANDD:   req_dcache_o.op = HPDCACHE_REQ_AMO_AND;
        AMO_ORW,AMO_ORD:     req_dcache_o.op = HPDCACHE_REQ_AMO_OR;
        AMO_MINW,AMO_MIND:   req_dcache_o.op = HPDCACHE_REQ_AMO_MIN;
        AMO_MAXW,AMO_MAXD:   req_dcache_o.op = HPDCACHE_REQ_AMO_MAX;
        AMO_MINWU,AMO_MINDU: req_dcache_o.op = HPDCACHE_REQ_AMO_MINU;
        AMO_MAXWU,AMO_MAXDU: req_dcache_o.op = HPDCACHE_REQ_AMO_MAXU;
        LD,LW,LWU,LH,LHU,LB,LBU,VLE,VLM,VL1R,VLEFF,VLSE,VLXE,FLD,FLW: req_dcache_o.op = HPDCACHE_REQ_LOAD;
        SD,SW,SH,SB,VSE,VSM,VS1R,FSW,FSD: req_dcache_o.op = HPDCACHE_REQ_STORE;
        default: req_dcache_o.op = HPDCACHE_REQ_LOAD;
    endcase
end

// Number of different sizes supported by the cache
localparam MAX_SIZES = $clog2(HPDCACHE_REQ_DATA_BYTES) + 1;

// CPU -> dCache data aligned to each size's natural alignment depending on the size & address
logic [HPDCACHE_REQ_DATA_WIDTH-1:0] aligned_data [MAX_SIZES-1:0];

generate
    for (genvar gv_size = 0; gv_size < MAX_SIZES; gv_size++) begin
        if (((1 << gv_size) * 8) <= riscv_pkg::VLEN) begin
            // If the requested size is smaller than the maximum generated by the core...
            if (((1 << gv_size) * 8) == HPDCACHE_REQ_DATA_WIDTH) begin
                // No shift needed, the request size is the whole request width's
                // and the core already aligns the data to the left, only select the bits used by gv_size
                assign aligned_data[gv_size] = req_cpu_dcache_i.data_rs2[(8 << gv_size)-1:0];
            end else begin
                // This will always be for smaller datatypes than HPDCACHE_REQ_DATA_WIDTH
                // because gv_size is generated for datatypes from byte to the whole request's width.
                // The following grabs only the bits used by gv_size (2^gv_size bytes)
                // and shifts it to align it to the request address and the size's align
                assign aligned_data[gv_size] =
                    req_cpu_dcache_i.data_rs2[(8 << gv_size)-1:0]
                        << {req_cpu_dcache_i.data_rs1[DCACHE_MAXELEM_LOG-1:gv_size], {{3+gv_size}{1'b0}}};
            end
        end else begin 
            // Else, if the requested size is larger than the maximum that the core can generate...
            // Send some dummy data. This, by construction, should never happen.
            // If you see these values in simulation or emulation... you f***** up.
            assign aligned_data[gv_size] = {{HPDCACHE_REQ_DATA_WIDTH/32}{32'hbadcab1e}};
        end
    end
endgenerate

// Select the write data depending on the request size
assign req_dcache_o.wdata = aligned_data[{req_cpu_dcache_i.mem_size[3], req_cpu_dcache_i.mem_size[1:0]}];

// *** Same as all of the above but for the byte enable signal ***

logic [HPDCACHE_REQ_DATA_BYTES-1:0] aligned_be [MAX_SIZES-1:0];

generate
    for (genvar gv_size = 0; gv_size < MAX_SIZES; gv_size++) begin
        if (((1 << gv_size) * 8) <= riscv_pkg::VLEN) begin
            // If the requested size is smaller than the maximum generated by the core...
            if (((1 << gv_size) * 8) == HPDCACHE_REQ_DATA_WIDTH) begin
                assign aligned_be[gv_size] = {{HPDCACHE_REQ_DATA_BYTES}{1'b1}};
            end else begin
                if (gv_size == 0) begin
                    assign aligned_be[gv_size] = {{1 << gv_size}{1'b1}} << {req_cpu_dcache_i.data_rs1[DCACHE_MAXELEM_LOG-1:gv_size]};
                end else begin
                    assign aligned_be[gv_size] =
                    {{1 << gv_size}{1'b1}} << {req_cpu_dcache_i.data_rs1[DCACHE_MAXELEM_LOG-1:gv_size], {{gv_size}{1'b0}}};
                end
            end
        end else begin 
            // If the requested size is larger than the maximum that the core
            // can generate, enable all bytes so that the mistake is obvious
            // during simulation/emulation (i.e. you can see the 0xbadcab1e).
            assign aligned_be[gv_size] = {{HPDCACHE_REQ_DATA_BYTES}{1'b1}};
        end
    end
endgenerate

assign req_dcache_o.be = aligned_be[{req_cpu_dcache_i.mem_size[3], req_cpu_dcache_i.mem_size[1:0]}];

assign req_dcache_o.addr_offset = req_cpu_dcache_i.data_rs1[(HPDCACHE_OFFSET_WIDTH+HPDCACHE_SET_WIDTH)-1:0],
       req_dcache_o.addr_tag = req_cpu_dcache_i.data_rs1[HPDCACHE_PA_WIDTH-1:(HPDCACHE_OFFSET_WIDTH+HPDCACHE_SET_WIDTH)];
// Request to HPDC. Pass only 2 bits as the sign extension process (see specs for LBU, LHU, LWU) is done in the mem_unit 
// HPDC does NOT extend the sign.
assign req_dcache_o.size = {req_cpu_dcache_i.mem_size[3], req_cpu_dcache_i.mem_size[1:0]}; // TODO: Core supports bigger memory sizes than HPDC!
assign req_dcache_o.sid = 3'b001;
assign req_dcache_o.tid = req_cpu_dcache_i.rd;
assign req_dcache_o.need_rsp = 1'b1;
assign req_dcache_o.phys_indexed = 1'b1;
assign req_dcache_o.pma.io = 1'b0;
assign req_dcache_o.pma.uncacheable = io_address_space;

// Unused signals on physically indexed requests
assign req_dcache_abort_o = 1'b0,
       req_dcache_tag_o = '0,
       req_dcache_pma_o = '0;

//-------------------------------------------------------------
// CPU Interface
//-------------------------------------------------------------

// Table holding the status of all the tags.
// This is a workaround to the HPDC not being able to process all the store
// requests the core is able to generate in time.
typedef enum logic {IDLE, PENDING} checker_state_t;
checker_state_t [127:0] transaction_table;


// Dcache interface to CPU 
assign resp_dcache_cpu_o.valid = dcache_valid_i;
assign resp_dcache_cpu_o.ready = dcache_ready_i & ~wait_resp_same_tag;
assign resp_dcache_cpu_o.io_address_space = io_address_space; // This should be done somewhere else...
assign resp_dcache_cpu_o.rd = rsp_dcache_i.tid;
assign resp_dcache_cpu_o.data = rsp_dcache_i.rdata;
assign resp_dcache_cpu_o.ordered = wbuf_empty_i;
// TODO: What about resp_dcache_cpu_o.error? Being tracked in issue #2.
// It's fine by now, the error signal is propagated from higher levels of the
// memory, which does *not* set it ever under any circumstance.

logic send, receive;

assign send    = core_req_valid_o && dcache_ready_i;
assign receive = dcache_valid_i;

//-PMU
assign dmem_is_store_o = (req_dcache_o.op == HPDCACHE_REQ_STORE) && send;
assign dmem_is_load_o  = (req_dcache_o.op == HPDCACHE_REQ_LOAD) && send;

`ifdef SIMULATION
logic [7:0] transactions_in_flight;
`endif

assign wait_resp_same_tag = transaction_table[req_dcache_o.tid] == PENDING;

always_ff @(posedge clk_i, negedge rstn_i) begin
    if (!rstn_i) begin
        for (int i = 0; i < 128; ++i) begin
            transaction_table[i] <= IDLE;
        end
        `ifdef SIMULATION
        transactions_in_flight <= 0;
        `endif
    end else begin
        if (send) begin
            `ifdef VERILATOR
            if (transaction_table[req_dcache_o.tid] == PENDING) begin
                $display("Transaction 0x%0h requested twice (time=%0t)", req_dcache_o.tid, $time);
                $fatal;
            end
            `endif

            transaction_table[req_dcache_o.tid] <= PENDING;
        end

        if (receive) begin
            `ifdef VERILATOR
            if (transaction_table[rsp_dcache_i.tid] == IDLE) begin
                $display("Transaction 0x%0h responded twice (time=%0t)", rsp_dcache_i.tid, $time);
                $fatal;
            end
            `endif

            transaction_table[rsp_dcache_i.tid] <= IDLE;
        end

        `ifdef SIMULATION
        transactions_in_flight <= transactions_in_flight + send - receive;
        `endif
    end
end

endmodule
//`default_nettype wire

