/*
 *  Authors       : Arnau Bigas
 *  Creation Date : July, 2023
 *  Description   : This file provides an AXI wrapper of the core, exposing the
 *                  memory hierarchy as a single AXI4 bus. Atomic operations are
 *                  implemented within this wrapper and thus needn't be
 *                  implemented upstream. This, however, implies that this
 *                  wrapper can only be used in single core applications.
 *                  Additionally, it also includes a bootrom.
 *  History      :
 */

import fpga_pkg::*, hpdcache_pkg::*;

module axi_wrapper (
    input logic clk_i,
    input logic rstn_i,

    AXI_BUS.Master axi_o,

    input logic time_irq_i,
    input logic [63:0] time_i
);

    // Bootrom wires
    logic [23:0] brom_req_address;
    logic brom_req_valid;
    logic brom_ready;
    logic [127:0] brom_resp_data;
    logic brom_resp_valid;

    // icache wires
    logic icache_l1_request_valid;
    logic icache_l2_response_valid;
    logic [drac_pkg::PHY_ADDR_SIZE-1:0] icache_l1_request_paddr;
    logic [511:0] icache_l2_response_data;

    logic core_icache_req_valid;
    logic core_icache_resp_valid;
    logic [drac_pkg::PHY_ADDR_SIZE-1:0] core_icache_request_paddr;
    logic [511:0] core_icache_response_data;
    logic [1:0] l2_response_seqnum;

    assign core_icache_response_data = brom_resp_valid ? brom_resp_data : icache_l2_response_data;
    assign core_icache_response_valid = brom_resp_valid | icache_l2_response_valid;
    assign icache_l1_request_paddr = core_icache_request_paddr;
    assign icache_l1_request_valid = core_icache_request_valid;

    //      Miss read interface
    logic                           mem_req_miss_read_ready;
    logic                           mem_req_miss_read_valid;
    sargantana_hpdc_pkg::hpdcache_mem_req_t    mem_req_miss_read;

    logic                           mem_resp_miss_read_ready;
    logic                           mem_resp_miss_read_valid;
    sargantana_hpdc_pkg::hpdcache_mem_resp_r_t mem_resp_miss_read;

    //      Write-buffer write interface
    logic                           mem_req_wbuf_write_ready;
    logic                           mem_req_wbuf_write_valid;
    sargantana_hpdc_pkg::hpdcache_mem_req_t    mem_req_wbuf_write;

    logic                           mem_req_wbuf_write_data_ready;
    logic                           mem_req_wbuf_write_data_valid;
    sargantana_hpdc_pkg::hpdcache_mem_req_w_t  mem_req_wbuf_write_data;

    logic                           mem_resp_wbuf_write_ready;
    logic                           mem_resp_wbuf_write_valid;
    sargantana_hpdc_pkg::hpdcache_mem_resp_w_t mem_resp_wbuf_write;

    //      Uncached read interface
    logic                           mem_req_uc_read_ready;
    logic                           mem_req_uc_read_valid;
    sargantana_hpdc_pkg::hpdcache_mem_req_t    mem_req_uc_read;
    sargantana_hpdc_pkg::hpdcache_mem_id_t     mem_req_uc_read_base_id;

    logic                           mem_resp_uc_read_ready;
    logic                           mem_resp_uc_read_valid;
    sargantana_hpdc_pkg::hpdcache_mem_resp_r_t mem_resp_uc_read;

    //      Uncached write interface
    logic                           mem_req_uc_write_ready;
    logic                           mem_req_uc_write_valid;
    sargantana_hpdc_pkg::hpdcache_mem_req_t    mem_req_uc_write;
    sargantana_hpdc_pkg::hpdcache_mem_id_t     mem_req_uc_write_base_id;

    logic                           mem_req_uc_write_data_ready;
    logic                           mem_req_uc_write_data_valid;
    sargantana_hpdc_pkg::hpdcache_mem_req_w_t  mem_req_uc_write_data;

    logic                           mem_resp_uc_write_ready;
    logic                           mem_resp_uc_write_valid;
    sargantana_hpdc_pkg::hpdcache_mem_resp_w_t mem_resp_uc_write;

    top_tile core_inst (
        .clk_i(clk_i),
        .rstn_i(rstn_i),
        .soft_rstn_i(rstn_i),
        .reset_addr_i(40'h0000000100),

        // Bootrom ports
        .brom_req_address_o(brom_req_address),
        .brom_req_valid_o(brom_req_valid),

        // icache ports
        .io_mem_acquire_valid(core_icache_request_valid),
        .io_mem_acquire_bits_addr_block(core_icache_request_paddr),
        .io_mem_grant_valid(core_icache_response_valid),
        .io_mem_grant_bits_data(core_icache_response_data),
        .io_mem_grant_bits_addr_beat(l2_response_seqnum),
        .io_mem_grant_inval(0),
        .io_mem_grant_inval_addr(0),

        // dmem ports

        // dMem miss-read interface
        .mem_req_miss_read_ready_i(mem_req_miss_read_ready),
        .mem_req_miss_read_valid_o(mem_req_miss_read_valid),
        .mem_req_miss_read_o(mem_req_miss_read),

        .mem_resp_miss_read_ready_o(mem_resp_miss_read_ready),
        .mem_resp_miss_read_valid_i(mem_resp_miss_read_valid),
        .mem_resp_miss_read_i(mem_resp_miss_read),

        // dMem writeback interface
        .mem_req_wbuf_write_ready_i(mem_req_wbuf_write_ready),
        .mem_req_wbuf_write_valid_o(mem_req_wbuf_write_valid),
        .mem_req_wbuf_write_o(mem_req_wbuf_write),

        .mem_req_wbuf_write_data_ready_i(mem_req_wbuf_write_data_ready),
        .mem_req_wbuf_write_data_valid_o(mem_req_wbuf_write_data_valid),
        .mem_req_wbuf_write_data_o(mem_req_wbuf_write_data),

        .mem_resp_wbuf_write_ready_o(mem_resp_wbuf_write_ready),
        .mem_resp_wbuf_write_valid_i(mem_resp_wbuf_write_valid),
        .mem_resp_wbuf_write_i(mem_resp_wbuf_write),

        // dMem uncacheable write interface
        .mem_req_uc_write_ready_i(mem_req_uc_write_ready),
        .mem_req_uc_write_valid_o(mem_req_uc_write_valid),
        .mem_req_uc_write_o(mem_req_uc_write),

        .mem_req_uc_write_data_ready_i(mem_req_uc_write_data_ready),
        .mem_req_uc_write_data_valid_o(mem_req_uc_write_data_valid),
        .mem_req_uc_write_data_o(mem_req_uc_write_data),

        .mem_resp_uc_write_ready_o(mem_resp_uc_write_ready),
        .mem_resp_uc_write_valid_i(mem_resp_uc_write_valid),
        .mem_resp_uc_write_i(mem_resp_uc_write),

        // dMem uncacheable read interface
        .mem_req_uc_read_ready_i(mem_req_uc_read_ready),
        .mem_req_uc_read_valid_o(mem_req_uc_read_valid),
        .mem_req_uc_read_o(mem_req_uc_read),

        .mem_resp_uc_read_ready_o(mem_resp_uc_read_ready),
        .mem_resp_uc_read_valid_i(mem_resp_uc_read_valid),
        .mem_resp_uc_read_i(mem_resp_uc_read),

        // Debug module
        .debug_contr_i('0),
        .debug_reg_i(¡0),
        .debug_contr_o(),
        .debug_reg_o(),

        .time_irq_i(time_irq_i),
        .irq_i(1'b0),
        .soft_irq_i(1'b0),
        .time_i(time_i)
    );

    bootrom brom(
        .clk(clk_i),
        .rstn(rstn_i),
        .brom_req_address_i(brom_req_address),
        .brom_req_valid_i(brom_req_valid),
        .brom_ready_o(brom_ready),
        .brom_resp_data_o(brom_resp_data),
        .brom_resp_valid_o(brom_resp_valid)
    );

    fpga_pkg::core_axi_req_t axi_req;
    fpga_pkg::core_axi_resp_t axi_resp;

    // Ojo! This breaks if hpdcache_pkg::HPDCACHE_MEM_TID_WIDTH <= (clog2(num_sets) + clog2(num_ways))!!!!
    assign mem_req_uc_read_base_id = '1;
    assign mem_req_uc_write_base_id = '1;

    axi_arbiter axi_arbiter_inst(
        .clk_i(clk_i),
        .rst_ni(rstn_i),

        // *** iCache ***

        .icache_miss_valid_i(icache_l1_request_valid),
        .icache_miss_paddr_i(icache_l1_request_paddr),
        .icache_miss_id_i(1 << (sargantana_hpdc_pkg::HPDCACHE_MEM_TID_WIDTH - 1)),

        .icache_miss_resp_valid_o(icache_l2_response_valid),
        .icache_miss_resp_data_o(icache_l2_response_data),
        .icache_miss_resp_beat_o(l2_response_seqnum),

        // *** dCache ***

        //      Miss-read interface
        .dcache_miss_ready_o(mem_req_miss_read_ready),
        .dcache_miss_valid_i(mem_req_miss_read_valid),
        .dcache_miss_i(mem_req_miss_read),

        .dcache_miss_resp_ready_i(mem_resp_miss_read_ready),
        .dcache_miss_resp_valid_o(mem_resp_miss_read_valid),
        .dcache_miss_resp_o(mem_resp_miss_read),

        //      Write-buffer write interface
        .dcache_wbuf_ready_o(mem_req_wbuf_write_ready),
        .dcache_wbuf_valid_i(mem_req_wbuf_write_valid),
        .dcache_wbuf_i(mem_req_wbuf_write),

        .dcache_wbuf_data_ready_o(mem_req_wbuf_write_data_ready),
        .dcache_wbuf_data_valid_i(mem_req_wbuf_write_data_valid),
        .dcache_wbuf_data_i(mem_req_wbuf_write_data),

        .dcache_wbuf_resp_ready_i(mem_resp_wbuf_write_ready),
        .dcache_wbuf_resp_valid_o(mem_resp_wbuf_write_valid),
        .dcache_wbuf_resp_o(mem_resp_wbuf_write),

        //      Uncached read interface
        .dcache_uc_read_ready_o(mem_req_uc_read_ready),
        .dcache_uc_read_valid_i(mem_req_uc_read_valid),
        .dcache_uc_read_i(mem_req_uc_read),
        .dcache_uc_read_id_i(mem_req_uc_read_base_id),

        .dcache_uc_read_resp_ready_i(mem_resp_uc_read_ready),
        .dcache_uc_read_resp_valid_o(mem_resp_uc_read_valid),
        .dcache_uc_read_resp_o(mem_resp_uc_read),

        //      Uncached write interface
        .dcache_uc_write_ready_o(mem_req_uc_write_ready),
        .dcache_uc_write_valid_i(mem_req_uc_write_valid),
        .dcache_uc_write_i(mem_req_uc_write),
        .dcache_uc_write_id_i(mem_req_uc_write_base_id),

        .dcache_uc_write_data_ready_o(mem_req_uc_write_data_ready),
        .dcache_uc_write_data_valid_i(mem_req_uc_write_data_valid),
        .dcache_uc_write_data_i(mem_req_uc_write_data),

        .dcache_uc_write_resp_ready_i(mem_resp_uc_write_ready),
        .dcache_uc_write_resp_valid_o(mem_resp_uc_write_valid),
        .dcache_uc_write_resp_o(mem_resp_uc_write),

        //  AXI port to upstream memory/peripherals
        .axi_req_o(axi_req),
        .axi_resp_i(axi_resp)
    );

    AXI_BUS #(
        .AXI_ADDR_WIDTH (64),
        .AXI_DATA_WIDTH (sargantana_hpdc_pkg::HPDCACHE_MEM_DATA_WIDTH),
        .AXI_ID_WIDTH   (sargantana_hpdc_pkg::HPDCACHE_MEM_TID_WIDTH),
        .AXI_USER_WIDTH (11)
    ) axi_core_to_atomic();

    `AXI_ASSIGN_FROM_REQ(axi_core_to_atomic, axi_req)
    `AXI_ASSIGN_TO_RESP(axi_resp, axi_core_to_atomic)

    AXI_BUS #(
        .AXI_ADDR_WIDTH (64),
        .AXI_DATA_WIDTH (sargantana_hpdc_pkg::HPDCACHE_MEM_DATA_WIDTH),
        .AXI_ID_WIDTH   (sargantana_hpdc_pkg::HPDCACHE_MEM_TID_WIDTH),
        .AXI_USER_WIDTH (11)
    ) axi_atomic_to_fpga();

    axi_riscv_atomics_wrap #(
        .AXI_ADDR_WIDTH(64),
        .AXI_DATA_WIDTH(sargantana_hpdc_pkg::HPDCACHE_MEM_DATA_WIDTH),
        .AXI_ID_WIDTH(sargantana_hpdc_pkg::HPDCACHE_MEM_TID_WIDTH),
        .AXI_USER_WIDTH(11),
        .AXI_MAX_READ_TXNS(1),
        .AXI_MAX_WRITE_TXNS(1),
        .RISCV_WORD_WIDTH(64)
    ) atomics_processor (
        .clk_i(clk_i),
        .rst_ni(rstn_i),
        .mst(axi_o),
        .slv(axi_core_to_atomic)
    );

endmodule
